package top_params_pkg;
    parameter NEW_FREQ_HZ     =           1;
    parameter DEFAULT_FREQ_HZ = 100_000_000;
    parameter WIDTH           =           3;
endpackage : top_params_pkg